module muladd1 inst(
	clk
	,a_0
	,a_1
	,a_2
	,a_3
	,b_0
	,b_1
	,b_2
	,b_3
	,sum

);


input clock;
input [15:0] a_0;
input [15:0] a_1;
input [15:0] a_2;
input [15:0] a_3;
input [15:0] b_0;
input [15:0] b_1;
input [15:0] b_2;
input [15:0] b_3;

output [15:0] sum;
























